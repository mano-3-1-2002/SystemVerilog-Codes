class transaction;
  rand bit [3:0]a;
  rand bit [3:0]b;
  bit [4:0]c;
endclass
