interface operation;
  logic [3:0]a;
  logic [3:0]b;
  logic [4:0]c;
endinterface
