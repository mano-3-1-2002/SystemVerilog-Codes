class transaction;
  rand bit d;
       bit clk;
  rand bit rst;
       bit q;
endclass
