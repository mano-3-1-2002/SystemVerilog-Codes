module add(input [3:0]a,[3:0]b,output[4:0] c);
  assign c = a+b;
endmodule
